library ieee;
use ieee.std_logic_1164.all;

entity multiplexer is
    port(
        i3  : in  std_logic_vector(31 downto 0);
        i2  : in  std_logic_vector(31 downto 0);
        i1  : in  std_logic_vector(31 downto 0);
        i0  : in  std_logic_vector(31 downto 0);
        sel : in  std_logic_vector(1 downto 0);
        o   : out std_logic_vector(31 downto 0)
    );
end multiplexer;

architecture synth of multiplexer is
begin

o <= i3 when sel = "00" else 
 	i2 when sel = "01" else
	i1 when sel = "10" else
	i0 when sel = "11";

end synth;
